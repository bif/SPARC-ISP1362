-------------------------------------------------------------------------------
-- Title      : Package Extension-Module
-- Project    : SCARTS - Scalable Processor for Embedded Applications in
--              Realtime Environment
-------------------------------------------------------------------------------
-- File       : pkg_display.vhd
-- Author     : Dipl. Ing. Martin Delvai
-- Company    : TU Wien - Institut fr Technische Informatik
-- Created    : 2002-02-11
-- Last update: 2011-10-20
-- Platform   : SUN Solaris
-------------------------------------------------------------------------------
-- Description:
-- Package for counter module
-------------------------------------------------------------------------------
-- Copyright (c) 2002 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2002-02-11  1.0      delvai	Created
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
-- LIBRARIES
-------------------------------------------------------------------------------

LIBRARY IEEE;
use IEEE.std_logic_1164.all;

use work.scarts_pkg.all;


-------------------------------------------------------------------------------
-- PACKAGE
-------------------------------------------------------------------------------

package pkg_counter is


-------------------------------------------------------------------------------
--                             CONSTANT
-------------------------------------------------------------------------------  

constant MY_CONFIGREG : natural := 3;
constant PRESCALER_REG : natural := 4;
constant CMD_COUNT : natural := 0;
constant CMD_CLEAR : natural := 1;

 
-------------------------------------------------------------------------------
-------------------------------------------------------------------------------
--                             COMPONENT
-------------------------------------------------------------------------------  
-------------------------------------------------------------------------------
    component ext_counter
      port (
        clk        : IN  std_logic;
        extsel     : in   std_ulogic;
        exti       : in  module_in_type;
        exto       : out module_out_type);
    end component;
  
   


end pkg_counter;
-------------------------------------------------------------------------------
--                             END PACKAGE
------------------------------------------------------------------------------- 
